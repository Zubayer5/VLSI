
interface Counter_Interface(input bit clk);
logic [15:0] data_in;
logic load;
logic enable;
logic up_down;
logic reset;
logic [15:0] data_out;
endinterface
