package memory_package;
`include"memory_stimulus.sv";
`include"memory_driver.sv";
`include"memory_monitor.sv";
`include"memory_agent.sv";
`include"memory_scoreboard.sv";
`include"memory_environment.sv";
`include"memory_test.sv";
endpackage
